library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity adder is
   port(A      : out std_logic;
        B      : out std_logic;
        C      : in  std_logic);
end adder;

architecture behv of adder is
   function rising_edge(c : in std_logic) return boolean;
begin
   process(A) is
   begin
      if A = B then
         if (not A) then
            C <= '0';
         end if;
      else
         C <= '1';
      end if;
   end process;
end behv;
